module ALU_testBench();
	wire [31:0]out;
	reg [31:0]inp1, inp2;
	reg [5:0]funct;
	
	
	// Calling module to test
	ALU alu(out, inp1, inp2, funct);
	
	
	
	// Test values
	initial begin
		inp1 = 32'b11111111111111111111111111111111; inp2 = 32'b00000000000000000000000000000000; funct = 6'b100000; #10;
		inp1 = 32'b11111111111111111111111111111100; inp2 = 32'b00000000000000000000000000000001; funct = 6'b100001; #10;
		inp1 = 32'b11111111111111111111111111111100; inp2 = 32'b11111111111111111111111111111000; funct = 6'b100010; #10;
		inp1 = 32'b10001111000011110000111100001111; inp2 = 32'b00111100001111000011110000111100; funct = 6'b100100; #10;
		inp1 = 32'b10001111000011110000111100001111; inp2 = 32'b00111100001111000011110000111100; funct = 6'b100101; #10;
		inp1 = 32'b10001111000011110000111100001111; inp2 = 32'b00111100001111000011110000111100; funct = 6'b101011; #10;
	end
	
	
	
	// Monitoring changes
	initial begin
		$monitor("Time=%2d, register0=%32b, register1=%32b, register2=%32b, funct=%6b", $time, inp1, inp2, out, funct);
	end
endmodule